///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: Flopenr (CLK=20)
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"

///////////////////////////////////////////////////////////////////////////////////
// Inputs: clk, reset, D, E (1-bit)
reg clk, reset, D, E;
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Output: Q (1-bit)
wire Q;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Component is CLOCKED
// Set clk period to 20 in wave
localparam CLK_PERIOD=20;
///////////////////////////////////////////////////////////////////////////////////

Flopenr myRegister(reset, clk, D, E, Q);

initial begin
/////////////////////////////////////////////////////////////////////////////
// Test: reset=1
$display("Testing reset: Q=0");
reset=1;  #(CLK_PERIOD/2);
verifyEqual(Q, 0);
/////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////
// Test: Falling edge
$display("Testing falling edge: Q=0");
reset=0;D=1;E=0; #(CLK_PERIOD/4);
verifyEqual(Q, 0);
/////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////
// Test: Enable off and rising edge
$display("Testing enable off with rising edge: Q=0");
#(CLK_PERIOD/2);
verifyEqual(Q, 0);
/////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////
// Test: Enable on and falling edge
$display("Testing enable on with falling edge: Q=0");
#(CLK_PERIOD/4);
E=1; #(CLK_PERIOD/4);
verifyEqual(Q, 0);
////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////
// Test: Enable on and rising edge
$display("Testing enable on with rising edge: Q=D");
#(CLK_PERIOD/2);
verifyEqual(Q, D);
/////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule

